----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:28:25 03/31/2013 
-- Design Name: 
-- Module Name:    main - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity main is
Port (
clk50 : in STD_LOGIC;
HS : out STD_LOGIC :='0';
VS : out STD_LOGIC :='0';

R : out  STD_LOGIC_VECTOR (2 downto 0);
G : out  STD_LOGIC_VECTOR (2 downto 0);
B : out  STD_LOGIC_VECTOR (1 downto 0);

xr : in STD_LOGIC :='0';
xl : in STD_LOGIC :='0';
yt : in STD_LOGIC :='0';
yb : in STD_LOGIC :='0';

SWITCH : in  STD_LOGIC_VECTOR (7 downto 0);

mplex: out STD_LOGIC_VECTOR (3 downto 0);
SEG : out std_logic_vector(6 downto 0));
end main;

architecture Behavioral of main is
signal Compteur_pixels: std_logic_vector(9 downto 0) :="0000000000";
signal Compteur_lignes: std_logic_vector(9 downto 0) :="0000000000";
signal origineX1: std_logic_vector(9 downto 0) :="0011001000";
signal origineY1: std_logic_vector(9 downto 0) :="0011001000";
signal origineX2: std_logic_vector(9 downto 0) :="0111110100";
signal origineY2: std_logic_vector(9 downto 0) :="0100101100";
signal Spot   :  std_logic_vector(8 downto 0) :="000000000";
signal color   :  std_logic_vector(8 downto 0) :="000000000";
signal tmp: std_logic_vector(3 downto 0) :="0000";
signal ds1:   std_logic_vector(3 downto 0):="0000";
signal us1:   std_logic_vector(3 downto 0):="0000";
signal ds2:   std_logic_vector(3 downto 0):="0000";
signal us2:   std_logic_vector(3 downto 0):="0000";
signal mp:   std_logic_vector(1 downto 0):="00";
signal score1: STD_LOGIC :='0';
signal score2: STD_LOGIC :='0';
signal time : std_logic_vector (25 downto 0):="00000000000000000000000000";
signal mtime: STD_LOGIC :='0';
signal timeout:   std_logic_vector(4 downto 0):="00000";
signal cpt: STD_LOGIC :='0';
signal Valide :  STD_LOGIC :='0';
signal clk25 :  STD_LOGIC :='0';
signal dpX :  STD_LOGIC :='0';
signal dpY :  STD_LOGIC :='0';
begin

--Clock 50Hz divis�e par 2 => 25Hz
process (clk50,clk25) 
begin
if clk50'event and clk50='1' then
	if clk25='1' then
		clk25<='0';
		else clk25<='1';
	end if;
	
	if score1='1' or score2='1' then
		timeout<="00000"; 
	end if;
	
	if (time = 49999999) then
		time<="00000000000000000000000000";
		timeout<=timeout+1;
		else
		time<=time+1;
	end if;
end if;
end process;

--Compteur pixels --Compteur lignes
process (clk25) 
begin
if clk25'event and clk25='1' then
	Compteur_pixels<= Compteur_pixels+1;
		if (Compteur_pixels= 799)then Compteur_pixels<= "0000000000"; 
		Compteur_lignes<= Compteur_lignes+1;
			if (Compteur_lignes= 519)then Compteur_lignes<= "0000000000";
			end if;
		end if;
end if;
end process;

--Affichage images
process (clk25)
CONSTANT tailleX :integer := 29;  
CONSTANT tailleY :integer := 29;
TYPE image is ARRAY(0 to tailleY, 0 to tailleX) OF std_logic_vector(8 downto 0);

CONSTANT chat : image :=(
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","111101111","100000000","111111111","111111111","111111111","111111111","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","110011110","100000000","011101111","010010110","010010110","010010101","001001101","011101111","100000000","110100110","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","010011110","001001101","001010110","010011110","010011110","010010110","001001101","010100110","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","111101111","010010110","010011111","010100111","011101111","010101111","010100111","010011111","001001101","010100101","111111111"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","011101111","010011110","010100111","011101111","011101111","011110111","011101111","010100111","010011110","001001100","111101110"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","011110111","001010110","001001110","001010110","010011110","010100111","011101111","011101111","010010110","001000100","101001101"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","111111111","011110111","001010101","001001101","001010110","010100111","010100111","010001101","001000100","011101111"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","111111111","100000000","100000000","110100110","001000100","001001101","010010110","010010101","010010101","001001101","011101110"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","101010101","001000011","001000011","010010101","010011110","010011111","001001100","101001100"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","111110111","100000000","100000000","100000000","100000000","111110111","010010101","001000100","010011110","010100111","010011110","001001100","001001011","111110110"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","111111111","100000000","100000000","111111111","011110111","111111111","100000000","010100110","001000100","010010101","010010101","001001100","000000011","001001011","111101110","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","010100110","110011101","100000000","111111111","100000000","011111111","010010110","001000100","000000011","000000010","010011101","001010101","001001100","010011110","001010110","001000101","010011110","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","110011101","101001100","111111111","010101110","001001100","000000100","010100110","001001101","001010100","010100110","001000100","001000011","001001100","010011110","001010101","000000010","000000011","001001101","001000100","001010100","011101110","111111111","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","110011101","001010101","001010110","010011110","010011101","000000010","000000011","001000100","000000011","001000100","001000011","001001100","010011111","010011110","010010101","010100110","010011110","001001100","001000100","101001100","111111111","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","110100110","010011111","010100101","001010110","000000011","001111111","001011101","000010100","001001011","000000011","001000011","010001101","010010101","011101111","010100110","010011110","011101111","010010101","001000011","010101110","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","111111111","100000000","110100111","010100111","011101110","010011111","001001100","001101110","001011101","010111111","000010100","000000011","001000100","010011110","010010101","010100110","011101111","010011110","010100111","010100111","001000011","001001100","100000000","111111111","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","011110111","010011110","010100110","011111111","010011111","010011110","001000100","001010101","001010100","001000100","001010110","001010110","001001101","001001100","010010110","011101111","010100110","010011110","010101111","001000100","000000011","111111111","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","011111111","001010101","001010110","011111111","010100110","010100111","001010101","001010101","010100111","010100111","010100111","010100110","010010110","000000011","010010101","010100111","010100111","010010101","010100111","001000011","000000010","011110111","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","111111111","101001101","010011110","001001101","011101111","011111111","010100110","010100111","010100110","010100110","010100111","011110110","011101111","001001101","001001100","010010101","010011110","010100111","010010101","010011111","001000011","000000010","011111111","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","110100111","001001100","010100111","010010110","001001100","011101111","011111111","011111111","011111111","011111111","011111111","011101111","001010110","001000011","001001101","010001101","010011110","010011110","001001101","001010101","000000001","001010100","100000000","111111111","100000000","100000000","100000000","100000000"),
("100000000","100000000","001001101","010001101","010001101","001000010","001010101","001001101","001010110","010100110","010100110","010100111","010010110","001001101","001001101","001000011","001001100","001001100","010011110","001010101","001000100","000000010","001001011","111101110","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","110011101","001001101","001000100","001000011","010011111","010011110","001000011","000000011","001000100","001000011","001001100","010011111","010011110","001001100","001000100","001000100","001010110","001000011","001001100","011101110","111111111","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","110011110","100000000","110011101","101001100","101010100","001001101","010010101","010010110","001000100","010011110","010001101","010001101","010001101","001001101","000000011","000000010","001000011","000000011","010011100","111110110","100000000","100000000","111111111","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","111111111","001001101","010010110","010001101","010011111","010011111","001001101","001000011","000000010","000000001","000000010","010011101","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","111111111","100000000","011101111","001001101","001000011","001001101","001001101","001010101","001010101","001010011","010100101","111111111","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","111111111","110011101","010100101","010011101","110010101","110101110","100000000","100000000","100000000","100000000","111110111","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000")
);

CONSTANT souris : image :=(
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100001001","100000000","100001001","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","001011011","101010010","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100001001","010100100","001010010","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","000001001","001010010","001010010","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100001001","000001001","001011011","010100100","001011011","000001001","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","001011011","001011011","001010010","010100100","010100100","001011011","010100100","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000001","001010011","001010011","001010011","001010010","001011011","010100100","001011011","010100100","010101101","010100100","010110110","001010010","000001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","001010011","010100110","010100110","010100110","001011100","010100100","010100100","010100100","010100100","011111111","010100100","001010010","001010010","001011011","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","001011101","010100110","010100110","010100110","010100110","001011100","010100100","010100100","010100100","001011100","001011100","001011100","001011100","001011011","101010010","100000000","101011011","100001001","100001001","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","001011100","010100110","010100110","001011101","001011100","001011011","010100011","010100100","001011011","000001001","001011100","001011100","001011100","001011011","100001001","010100100","010101101","010100100","001011011","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","001010011","010101110","010100110","001011100","010100100","010100100","010100100","010100100","001011011","000001001","000000000","000000000","001011100","001010010","010101101","010101101","001011011","001011011","101010010","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","001011100","010100110","010100101","010101101","011110110","010101101","001011011","010100101","001011101","000001110","000001011","001011100","010101101","011110110","101011011","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100001001","100000000","100001010","001011100","001011100","010100100","010100100","010101101","010101101","010100100","001011100","001010101","000001100","010100100","010101101","010101101","100001001","100000000","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","101011101","100000000","100000001","100001010","101010011","101010010","001011011","010101101","011110110","010101110","010100100","010100100","010100101","001100100","101010010","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","101011011","010101101","011110110","011110110","010101110","010101111","010101111","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100001001","100001001","100001001","100001010","001010010","101010011","100000000","001010010","010101101","011110110","010101111","010110111","010101110","001011011","001011011","001010011","100001010","100001010","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","101010011","100000000","100000001","100001001","100001010","100001010","001010011","001010011","010100100","011110110","010101110","010110111","010110111","010101110","010100100","010100101","010100101","001011101","100001010","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100001001","100001001","010101101","011110110","010110110","010101111","010110111","010110111","010100101","001011100","010100110","010100110","101010011","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100001001","001011011","010101101","010100100","011110110","010110110","010101111","010110111","010110111","001100101","001011011","001011100","010100110","001011100","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","101011011","010101101","010101101","010110110","011110110","010101110","010110111","010110111","001100101","101010010","100001001","001011100","001011101","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","101011011","010101101","010100100","011110110","011110110","010101101","001011011","000010010","100000000","100000000","100000000","100001001","100000001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","101010010","001010010","010101101","010100100","101011011","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100001001","101010010","100001001","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000"),
("100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000","100000000")
);
variable Ligne1:integer:=0;
variable Ligne2:integer:=0;
variable Pixel1:integer:=0;
variable Pixel2:integer:=0;

begin
if clk25'event and clk25='1' then
		if Compteur_pixels >= origineX1 and compteur_pixels < origineX1 +tailleX and compteur_lignes >= origineY1
		 and compteur_lignes < origineY1 + tailleY  then
			if chat(ligne1,Pixel1)(8)='1' then
			Spot <= color;
			else
			Spot <= chat (ligne1,Pixel1);
			end if;
			Pixel1 := Pixel1+1;
			if pixel1 = tailleX then pixel1 := 0; ligne1 := ligne1 + 1;
					if ligne1 = tailleY then ligne1 := 0;
					end if;
				end if;
			elsif Compteur_pixels >= origineX2 and compteur_pixels < origineX2 +tailleX and compteur_lignes >= origineY2
			and compteur_lignes < origineY2 + tailleY  then
				if souris(ligne2,Pixel2)(8)='1' then
				Spot <= color;
				else
				Spot <= souris (ligne2,Pixel2);
				end if;
			Pixel2 := Pixel2+1;
			if pixel2 = tailleX then pixel2 := 0; ligne2 := ligne2 + 1;
					if ligne2 = tailleY then ligne2 := 0;
					end if;
				end if;
			else 
			Spot <= color;
		end if;
		
		--D�placement � la fin de l'affichage
		if Compteur_lignes= 519 and Compteur_pixels= 799 then
			--D�placement chat
			if origineX1 + tailleX + 1 <783 and xr='1' then origineX1 <= origineX1 +1; --Mouvement X1
			end if;
			if origineX1 >144 and xl='1' then origineX1 <= origineX1 -1;
			end if;
			
			if origineY1 + tailleY + 1 <510 and yb='1' then origineY1 <= origineY1 +1; --Mouvement Y1
			end if;
			if origineY1 >31 and yt='1' then origineY1 <= origineY1 -1;
			end if;
			
			--D�placement souris
			if origineX2 + tailleX + 1 >783 then dpX<='1'; --Mouvement X2
			end if;
			if origineX2 <144 then dpX<='0';
			end if;
			
			if dpX='0' then origineX2 <= origineX2 +1;
			else origineX2 <= origineX2 -1;
			end if;
			
			if origineY2 + tailleY + 1 >510 then dpY<='1'; --Mouvement Y2
			end if;
			if origineY2 <31 then dpY<='0';
			end if;
			
			if dpY='0' then origineY2 <= origineY2 +1;
			else origineY2 <= origineY2 -1;
			end if;
		end if;
		score1<='0';
		score2<='0';
		--Le chat mange la souris
		if origineX1+tailleX>origineX2 and origineX1-tailleX<origineX2 
		and origineY1+tailleY>origineY2 and origineY1-tailleY<origineY2 then
			origineX1  <="0011001000";
			origineY1 <="0011001000";
			origineX2 <="0111110100";
			origineY2 <="0100101100";
			score1<='1';
		end if;
		
		--La souris gagne temps>30 sec
		if timeout=30 then
		origineX1  <="0011001000";
		origineY1 <="0011001000";
		origineX2 <="0111110100";
		origineY2 <="0100101100";
		score2<='1';
		end if;
end if;
end process;

mtime<=time(15);
process(clk25)
 	begin
		if mtime'event and mtime='1' then
		mp<=mp+1;
		end if;
end process;

--Compteur score
process(clk25)
 	begin
		if clk25'event and clk25='1' then
		if score1='1' then
		us1<=us1+1;
		end if;
		if score2='1' then
		us2<=us2+1;
		end if;
			if (us1=9) then 
			ds1<=ds1+1;
			us1 <= "0000";
				if (ds1=9) then
				ds1 <= "0000";
				end if;
			end if;
			if (us2=9) then
			ds2<=ds2+1;
			us2 <= "0000";
				if (ds2=9) then
				ds2 <= "0000";
				end if;
			end if;
		end if;
end process;
		 	 
		with mp select			
		mplex <= "1110" when "00",
		"1101" when "01",
		"1011" when "10",
		"0111" when "11",
		"1111" when others;	
	
	   with mp select
		tmp <= us1 when "00",
		ds1 when "01",
		us2 when "10",
		ds2 when "11",
		"0000" when others;
	     
	--Affichage couleur
	Valide <= '1' when (Compteur_pixels>=144 and Compteur_pixels<783 and Compteur_lignes>=31 and Compteur_lignes<510) else '0';
	HS <= '0' when Compteur_pixels < 96 else '1';
	VS <= '0' when Compteur_lignes < 2 else '1';
	R(0) <= '1' when (Valide='1' and  Spot(0)='1') else '0';
	R(1) <= '1' when (Valide='1' and  Spot(1)='1') else '0';
	R(2) <= '1' when (Valide='1' and  Spot(2)='1') else '0';
	G(0) <= '1' when (Valide='1' and  Spot(3)='1') else '0';
	G(1) <= '1' when (Valide='1' and  Spot(4)='1') else '0';
	G(2) <= '1' when (Valide='1' and  Spot(5)='1') else '0';
	B(0) <= '1' when (Valide='1' and  Spot(6)='1') else '0';
	B(1) <= '1' when (Valide='1' and  Spot(7)='1') else '0';
	
	--Choix couleur de fond
	color(0)<='1' when SWITCH(0)='1' else '0';
	color(1)<='1' when SWITCH(1)='1' else '0';
	color(2)<='1' when SWITCH(2)='1' else '0';
	color(3)<='1' when SWITCH(3)='1' else '0';
	color(4)<='1' when SWITCH(4)='1' else '0';
	color(5)<='1' when SWITCH(5)='1' else '0';
	color(6)<='1' when SWITCH(6)='1' else '0';
	color(7)<='1' when SWITCH(7)='1' else '0';

  SEG<="1000000" when tmp ="0000"
		else "1111001" when tmp ="0001"
		else "0100100"	when tmp ="0010"
		else "0110000"	when tmp ="0011"
		else "0011001"	when tmp ="0100"
		else "0010010" when tmp ="0101"
		else "0000010"	when tmp ="0110"
		else "1111000" when tmp ="0111"
		else "0000000" when tmp ="1000"
		else "0010000"	when tmp ="1001"
		else "0111111";
		

end Behavioral;